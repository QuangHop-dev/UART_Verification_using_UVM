package UART_pkg;
    import uvm_pkg::*;
    
    `include "uvm_macros.svh"

    `include "sequence_item.sv"
    `include "sequence.sv"
    `include "sequencer.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "coverage_collector.sv"
    `include "scoreboard.sv"
    `include "agent.sv"
    `include "env.sv"
    `include "test.sv"
	
endpackage: UART_pkg
